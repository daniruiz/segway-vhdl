

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity control_motores is
    generic ( n_bits_datos : integer := 8 );
    port    ( reloj        : in std_logic;
              x_gyro       : in std_logic_vector (n_bits_datos-1 downto 0); -- inclinación
              y_gyro       : in std_logic_vector (n_bits_datos-1 downto 0); -- giro
              y_accel      : in std_logic_vector (n_bits_datos-1 downto 0);
              z_accel      : in std_logic_vector (n_bits_datos-1 downto 0);
              velocidad_a  : out std_logic_vector (7 downto 0);
              l298n_in1    : out std_logic; -- sentido motor a _0
              l298n_in2    : out std_logic; -- sentido motor a _1
              l298n_in3    : out std_logic; -- sentido motor b _0
              l298n_in4    : out std_logic; -- sentido motor b _1
              velocidad_b  : out std_logic_vector (7 downto 0);
              
              kpUp         : in std_logic;
              kdUP         : in std_logic;
              kiUP         : in std_logic;
              
              KP           : inout integer;
              KD           : inout integer;
              KI           : inout integer );
end control_motores;

architecture comportamiento of control_motores is

    constant decimales         : integer   := 1000;
    constant timeChange        : integer   := 1; -- 0.1 ns
    constant vel_offset        : integer   := 70;
    constant gyro_gain         : integer   := 91; -- (65 * 127 * 2 / 180);
    constant A                 : integer   := 987;
    constant dt                : integer   := 10; -- 10 ms => 10/1000 s
 
    signal velocidad_a_integer : integer;
    signal velocidad_b_integer : integer;

    function calc_angulo_crudo (y_accel : integer; z_accel : integer) return integer is
        type t_valores is array(0 to 10000) of integer;
        -- 180_deg := 127*2;
        -- atan( y_accel / z_accel ) / pi * 180_deg;   *1000 para 3 decimales
        variable valores : t_valores := (0,808,1616,2424,3232,4039,4845,5650,6454,7257,8058,8857,9655,10451,11246,12037,12827,13614,14398,15180,15959,16735,17508,18277,19043,19806,20565,21321,22072,22820,23564,24304,25039,25770,26497,27220,27938,28651,29360,30064,30764,31458,32148,32833,33513,34188,34857,35522,36182,36836,37486,38130,38769,39403,40031,40655,41273,41886,42493,43096,43693,44285,44871,45453,46029,46600,47166,47726,48282,48832,49377,49917,50452,50982,51507,52027,52542,53052,53557,54057,54553,55043,55529,56010,56487,56958,57425,57888,58346,58799,59248,59693,60133,60568,61000,61427,61850,62268,62683,63093,63500,63902,64300,64694,65085,65471,65854,66233,66608,66979,67347,67711,68071,68428,68781,69131,69478,69821,70160,70496,70829,71159,71486,71809,72129,72446,72760,73071,73379,73684,73986,74285,74581,74875,75165,75453,75738,76021,76300,76577,76852,77124,77393,77660,77924,78186,78445,78702,78957,79209,79459,79707,79952,80195,80436,80675,80911,81146,81378,81608,81836,82062,82287,82509,82729,82947,83163,83377,83590,83800,84009,84216,84421,84625,84826,85026,85224,85421,85616,85809,86000,86190,86378,86565,86750,86934,87116,87296,87475,87653,87829,88004,88177,88349,88519,88688,88856,89022,89187,89351,89513,89674,89834,89993,90150,90306,90461,90614,90767,90918,91068,91217,91364,91511,91657,91801,91944,92086,92227,92367,92506,92644,92781,92917,93052,93186,93319,93451,93581,93711,93840,93968,94096,94222,94347,94472,94595,94718,94839,94960,95080,95200,95318,95435,95552,95668,95783,95897,96011,96123,96235,96346,96457,96566,96675,96783,96891,96997,97103,97209,97313,97417,97520,97623,97724,97826,97926,98026,98125,98223,98321,98419,98515,98611,98706,98801,98895,98989,99082,99174,99266,99357,99448,99538,99627,99716,99804,99892,99979,100066,100152,100238,100323,100408,100492,100575,100658,100741,100823,100905,100986,101066,101146,101226,101305,101384,101462,101540,101617,101694,101771,101847,101922,101997,102072,102146,102220,102293,102366,102439,102511,102583,102654,102725,102796,102866,102935,103005,103074,103142,103210,103278,103346,103413,103479,103546,103612,103677,103743,103807,103872,103936,104000,104064,104127,104190,104252,104314,104376,104438,104499,104560,104620,104680,104740,104800,104859,104918,104977,105035,105093,105151,105208,105266,105323,105379,105435,105491,105547,105603,105658,105713,105767,105822,105876,105930,105983,106036,106089,106142,106195,106247,106299,106351,106402,106453,106504,106555,106606,106656,106706,106756,106805,106854,106903,106952,107001,107049,107097,107145,107193,107240,107287,107334,107381,107428,107474,107520,107566,107612,107657,107703,107748,107793,107837,107882,107926,107970,108014,108058,108101,108144,108188,108230,108273,108316,108358,108400,108442,108484,108525,108567,108608,108649,108690,108731,108771,108811,108851,108891,108931,108971,109010,109050,109089,109128,109166,109205,109244,109282,109320,109358,109396,109433,109471,109508,109545,109582,109619,109656,109693,109729,109765,109801,109837,109873,109909,109944,109980,110015,110050,110085,110120,110154,110189,110223,110258,110292,110326,110359,110393,110427,110460,110493,110527,110560,110593,110625,110658,110690,110723,110755,110787,110819,110851,110883,110915,110946,110977,111009,111040,111071,111102,111133,111163,111194,111224,111255,111285,111315,111345,111375,111405,111434,111464,111493,111523,111552,111581,111610,111639,111668,111696,111725,111753,111782,111810,111838,111866,111894,111922,111950,111977,112005,112032,112060,112087,112114,112141,112168,112195,112222,112248,112275,112301,112328,112354,112380,112406,112432,112458,112484,112510,112535,112561,112586,112612,112637,112662,112687,112712,112737,112762,112787,112812,112836,112861,112885,112910,112934,112958,112982,113006,113030,113054,113078,113101,113125,113149,113172,113195,113219,113242,113265,113288,113311,113334,113357,113380,113402,113425,113448,113470,113492,113515,113537,113559,113581,113603,113625,113647,113669,113691,113712,113734,113755,113777,113798,113820,113841,113862,113883,113904,113925,113946,113967,113988,114009,114029,114050,114070,114091,114111,114132,114152,114172,114192,114212,114232,114252,114272,114292,114312,114332,114351,114371,114390,114410,114429,114449,114468,114487,114506,114525,114545,114564,114582,114601,114620,114639,114658,114676,114695,114714,114732,114750,114769,114787,114805,114824,114842,114860,114878,114896,114914,114932,114950,114968,114985,115003,115021,115038,115056,115073,115091,115108,115125,115143,115160,115177,115194,115211,115228,115245,115262,115279,115296,115313,115330,115346,115363,115380,115396,115413,115429,115446,115462,115478,115495,115511,115527,115543,115559,115575,115591,115607,115623,115639,115655,115671,115686,115702,115718,115733,115749,115765,115780,115796,115811,115826,115842,115857,115872,115887,115902,115918,115933,115948,115963,115978,115993,116007,116022,116037,116052,116067,116081,116096,116110,116125,116140,116154,116168,116183,116197,116212,116226,116240,116254,116268,116283,116297,116311,116325,116339,116353,116367,116381,116394,116408,116422,116436,116449,116463,116477,116490,116504,116517,116531,116544,116558,116571,116585,116598,116611,116624,116638,116651,116664,116677,116690,116703,116716,116729,116742,116755,116768,116781,116794,116807,116819,116832,116845,116857,116870,116883,116895,116908,116920,116933,116945,116958,116970,116982,116995,117007,117019,117032,117044,117056,117068,117080,117092,117104,117117,117129,117140,117152,117164,117176,117188,117200,117212,117224,117235,117247,117259,117270,117282,117294,117305,117317,117328,117340,117351,117363,117374,117385,117397,117408,117420,117431,117442,117453,117464,117476,117487,117498,117509,117520,117531,117542,117553,117564,117575,117586,117597,117608,117619,117629,117640,117651,117662,117673,117683,117694,117705,117715,117726,117736,117747,117757,117768,117778,117789,117799,117810,117820,117831,117841,117851,117861,117872,117882,117892,117902,117913,117923,117933,117943,117953,117963,117973,117983,117993,118003,118013,118023,118033,118043,118053,118063,118072,118082,118092,118102,118112,118121,118131,118141,118150,118160,118170,118179,118189,118198,118208,118217,118227,118236,118246,118255,118265,118274,118283,118293,118302,118311,118321,118330,118339,118348,118358,118367,118376,118385,118394,118403,118412,118422,118431,118440,118449,118458,118467,118476,118485,118493,118502,118511,118520,118529,118538,118547,118555,118564,118573,118582,118590,118599,118608,118616,118625,118634,118642,118651,118660,118668,118677,118685,118694,118702,118711,118719,118728,118736,118744,118753,118761,118770,118778,118786,118795,118803,118811,118819,118828,118836,118844,118852,118860,118869,118877,118885,118893,118901,118909,118917,118925,118933,118941,118949,118957,118965,118973,118981,118989,118997,119005,119013,119020,119028,119036,119044,119052,119060,119067,119075,119083,119091,119098,119106,119114,119121,119129,119137,119144,119152,119159,119167,119174,119182,119190,119197,119205,119212,119219,119227,119234,119242,119249,119257,119264,119271,119279,119286,119293,119301,119308,119315,119323,119330,119337,119344,119352,119359,119366,119373,119380,119387,119395,119402,119409,119416,119423,119430,119437,119444,119451,119458,119465,119472,119479,119486,119493,119500,119507,119514,119521,119528,119535,119541,119548,119555,119562,119569,119576,119582,119589,119596,119603,119609,119616,119623,119630,119636,119643,119650,119656,119663,119670,119676,119683,119689,119696,119703,119709,119716,119722,119729,119735,119742,119748,119755,119761,119768,119774,119781,119787,119793,119800,119806,119813,119819,119825,119832,119838,119844,119851,119857,119863,119869,119876,119882,119888,119894,119901,119907,119913,119919,119925,119932,119938,119944,119950,119956,119962,119968,119974,119981,119987,119993,119999,120005,120011,120017,120023,120029,120035,120041,120047,120053,120059,120065,120071,120076,120082,120088,120094,120100,120106,120112,120118,120123,120129,120135,120141,120147,120153,120158,120164,120170,120176,120181,120187,120193,120198,120204,120210,120216,120221,120227,120233,120238,120244,120249,120255,120261,120266,120272,120277,120283,120289,120294,120300,120305,120311,120316,120322,120327,120333,120338,120344,120349,120355,120360,120366,120371,120376,120382,120387,120393,120398,120403,120409,120414,120419,120425,120430,120435,120441,120446,120451,120457,120462,120467,120472,120478,120483,120488,120493,120499,120504,120509,120514,120519,120525,120530,120535,120540,120545,120550,120555,120561,120566,120571,120576,120581,120586,120591,120596,120601,120606,120611,120616,120621,120626,120631,120636,120641,120646,120651,120656,120661,120666,120671,120676,120681,120686,120691,120696,120701,120706,120711,120715,120720,120725,120730,120735,120740,120745,120749,120754,120759,120764,120769,120773,120778,120783,120788,120792,120797,120802,120807,120811,120816,120821,120826,120830,120835,120840,120844,120849,120854,120858,120863,120868,120872,120877,120882,120886,120891,120895,120900,120905,120909,120914,120918,120923,120927,120932,120936,120941,120946,120950,120955,120959,120964,120968,120973,120977,120982,120986,120990,120995,120999,121004,121008,121013,121017,121021,121026,121030,121035,121039,121043,121048,121052,121057,121061,121065,121070,121074,121078,121083,121087,121091,121096,121100,121104,121108,121113,121117,121121,121126,121130,121134,121138,121143,121147,121151,121155,121159,121164,121168,121172,121176,121180,121185,121189,121193,121197,121201,121205,121210,121214,121218,121222,121226,121230,121234,121238,121242,121247,121251,121255,121259,121263,121267,121271,121275,121279,121283,121287,121291,121295,121299,121303,121307,121311,121315,121319,121323,121327,121331,121335,121339,121343,121347,121351,121355,121359,121363,121367,121370,121374,121378,121382,121386,121390,121394,121398,121402,121405,121409,121413,121417,121421,121425,121429,121432,121436,121440,121444,121448,121451,121455,121459,121463,121467,121470,121474,121478,121482,121485,121489,121493,121497,121500,121504,121508,121512,121515,121519,121523,121526,121530,121534,121538,121541,121545,121549,121552,121556,121560,121563,121567,121571,121574,121578,121581,121585,121589,121592,121596,121599,121603,121607,121610,121614,121617,121621,121625,121628,121632,121635,121639,121642,121646,121649,121653,121656,121660,121664,121667,121671,121674,121678,121681,121685,121688,121692,121695,121698,121702,121705,121709,121712,121716,121719,121723,121726,121730,121733,121736,121740,121743,121747,121750,121753,121757,121760,121764,121767,121770,121774,121777,121780,121784,121787,121791,121794,121797,121801,121804,121807,121811,121814,121817,121821,121824,121827,121830,121834,121837,121840,121844,121847,121850,121853,121857,121860,121863,121867,121870,121873,121876,121879,121883,121886,121889,121892,121896,121899,121902,121905,121908,121912,121915,121918,121921,121924,121928,121931,121934,121937,121940,121943,121947,121950,121953,121956,121959,121962,121965,121969,121972,121975,121978,121981,121984,121987,121990,121993,121997,122000,122003,122006,122009,122012,122015,122018,122021,122024,122027,122030,122033,122036,122039,122043,122046,122049,122052,122055,122058,122061,122064,122067,122070,122073,122076,122079,122082,122085,122088,122091,122094,122097,122100,122102,122105,122108,122111,122114,122117,122120,122123,122126,122129,122132,122135,122138,122141,122144,122147,122149,122152,122155,122158,122161,122164,122167,122170,122173,122175,122178,122181,122184,122187,122190,122193,122195,122198,122201,122204,122207,122210,122213,122215,122218,122221,122224,122227,122229,122232,122235,122238,122241,122243,122246,122249,122252,122255,122257,122260,122263,122266,122268,122271,122274,122277,122280,122282,122285,122288,122291,122293,122296,122299,122301,122304,122307,122310,122312,122315,122318,122320,122323,122326,122329,122331,122334,122337,122339,122342,122345,122347,122350,122353,122355,122358,122361,122363,122366,122369,122371,122374,122377,122379,122382,122384,122387,122390,122392,122395,122398,122400,122403,122405,122408,122411,122413,122416,122418,122421,122424,122426,122429,122431,122434,122437,122439,122442,122444,122447,122449,122452,122454,122457,122460,122462,122465,122467,122470,122472,122475,122477,122480,122482,122485,122487,122490,122492,122495,122497,122500,122502,122505,122507,122510,122512,122515,122517,122520,122522,122525,122527,122530,122532,122535,122537,122540,122542,122545,122547,122549,122552,122554,122557,122559,122562,122564,122566,122569,122571,122574,122576,122579,122581,122583,122586,122588,122591,122593,122595,122598,122600,122603,122605,122607,122610,122612,122615,122617,122619,122622,122624,122626,122629,122631,122633,122636,122638,122640,122643,122645,122648,122650,122652,122655,122657,122659,122662,122664,122666,122668,122671,122673,122675,122678,122680,122682,122685,122687,122689,122692,122694,122696,122698,122701,122703,122705,122708,122710,122712,122714,122717,122719,122721,122723,122726,122728,122730,122732,122735,122737,122739,122741,122744,122746,122748,122750,122753,122755,122757,122759,122761,122764,122766,122768,122770,122773,122775,122777,122779,122781,122784,122786,122788,122790,122792,122795,122797,122799,122801,122803,122805,122808,122810,122812,122814,122816,122818,122821,122823,122825,122827,122829,122831,122833,122836,122838,122840,122842,122844,122846,122848,122851,122853,122855,122857,122859,122861,122863,122865,122868,122870,122872,122874,122876,122878,122880,122882,122884,122886,122889,122891,122893,122895,122897,122899,122901,122903,122905,122907,122909,122911,122913,122915,122918,122920,122922,122924,122926,122928,122930,122932,122934,122936,122938,122940,122942,122944,122946,122948,122950,122952,122954,122956,122958,122960,122962,122964,122966,122968,122970,122972,122974,122976,122978,122980,122982,122984,122986,122988,122990,122992,122994,122996,122998,123000,123002,123004,123006,123008,123010,123012,123014,123016,123018,123020,123022,123024,123026,123028,123030,123032,123034,123036,123037,123039,123041,123043,123045,123047,123049,123051,123053,123055,123057,123059,123061,123063,123064,123066,123068,123070,123072,123074,123076,123078,123080,123082,123083,123085,123087,123089,123091,123093,123095,123097,123099,123100,123102,123104,123106,123108,123110,123112,123114,123115,123117,123119,123121,123123,123125,123127,123128,123130,123132,123134,123136,123138,123140,123141,123143,123145,123147,123149,123151,123152,123154,123156,123158,123160,123161,123163,123165,123167,123169,123171,123172,123174,123176,123178,123180,123181,123183,123185,123187,123189,123190,123192,123194,123196,123198,123199,123201,123203,123205,123206,123208,123210,123212,123214,123215,123217,123219,123221,123222,123224,123226,123228,123229,123231,123233,123235,123236,123238,123240,123242,123243,123245,123247,123249,123250,123252,123254,123256,123257,123259,123261,123263,123264,123266,123268,123269,123271,123273,123275,123276,123278,123280,123281,123283,123285,123287,123288,123290,123292,123293,123295,123297,123298,123300,123302,123304,123305,123307,123309,123310,123312,123314,123315,123317,123319,123320,123322,123324,123325,123327,123329,123330,123332,123334,123335,123337,123339,123340,123342,123344,123345,123347,123349,123350,123352,123353,123355,123357,123358,123360,123362,123363,123365,123367,123368,123370,123371,123373,123375,123376,123378,123380,123381,123383,123384,123386,123388,123389,123391,123392,123394,123396,123397,123399,123401,123402,123404,123405,123407,123408,123410,123412,123413,123415,123416,123418,123420,123421,123423,123424,123426,123428,123429,123431,123432,123434,123435,123437,123439,123440,123442,123443,123445,123446,123448,123449,123451,123453,123454,123456,123457,123459,123460,123462,123463,123465,123467,123468,123470,123471,123473,123474,123476,123477,123479,123480,123482,123483,123485,123486,123488,123490,123491,123493,123494,123496,123497,123499,123500,123502,123503,123505,123506,123508,123509,123511,123512,123514,123515,123517,123518,123520,123521,123523,123524,123526,123527,123529,123530,123532,123533,123535,123536,123538,123539,123541,123542,123543,123545,123546,123548,123549,123551,123552,123554,123555,123557,123558,123560,123561,123563,123564,123565,123567,123568,123570,123571,123573,123574,123576,123577,123579,123580,123581,123583,123584,123586,123587,123589,123590,123592,123593,123594,123596,123597,123599,123600,123602,123603,123604,123606,123607,123609,123610,123612,123613,123614,123616,123617,123619,123620,123621,123623,123624,123626,123627,123628,123630,123631,123633,123634,123635,123637,123638,123640,123641,123642,123644,123645,123647,123648,123649,123651,123652,123654,123655,123656,123658,123659,123660,123662,123663,123665,123666,123667,123669,123670,123671,123673,123674,123676,123677,123678,123680,123681,123682,123684,123685,123686,123688,123689,123691,123692,123693,123695,123696,123697,123699,123700,123701,123703,123704,123705,123707,123708,123709,123711,123712,123713,123715,123716,123717,123719,123720,123721,123723,123724,123725,123727,123728,123729,123731,123732,123733,123735,123736,123737,123739,123740,123741,123742,123744,123745,123746,123748,123749,123750,123752,123753,123754,123756,123757,123758,123759,123761,123762,123763,123765,123766,123767,123768,123770,123771,123772,123774,123775,123776,123777,123779,123780,123781,123783,123784,123785,123786,123788,123789,123790,123792,123793,123794,123795,123797,123798,123799,123800,123802,123803,123804,123805,123807,123808,123809,123811,123812,123813,123814,123816,123817,123818,123819,123821,123822,123823,123824,123826,123827,123828,123829,123831,123832,123833,123834,123835,123837,123838,123839,123840,123842,123843,123844,123845,123847,123848,123849,123850,123851,123853,123854,123855,123856,123858,123859,123860,123861,123862,123864,123865,123866,123867,123869,123870,123871,123872,123873,123875,123876,123877,123878,123879,123881,123882,123883,123884,123885,123887,123888,123889,123890,123891,123893,123894,123895,123896,123897,123899,123900,123901,123902,123903,123904,123906,123907,123908,123909,123910,123912,123913,123914,123915,123916,123917,123919,123920,123921,123922,123923,123924,123926,123927,123928,123929,123930,123931,123933,123934,123935,123936,123937,123938,123940,123941,123942,123943,123944,123945,123947,123948,123949,123950,123951,123952,123953,123955,123956,123957,123958,123959,123960,123961,123963,123964,123965,123966,123967,123968,123969,123971,123972,123973,123974,123975,123976,123977,123978,123980,123981,123982,123983,123984,123985,123986,123987,123989,123990,123991,123992,123993,123994,123995,123996,123998,123999,124000,124001,124002,124003,124004,124005,124006,124008,124009,124010,124011,124012,124013,124014,124015,124016,124017,124019,124020,124021,124022,124023,124024,124025,124026,124027,124028,124029,124031,124032,124033,124034,124035,124036,124037,124038,124039,124040,124041,124043,124044,124045,124046,124047,124048,124049,124050,124051,124052,124053,124054,124055,124056,124058,124059,124060,124061,124062,124063,124064,124065,124066,124067,124068,124069,124070,124071,124072,124074,124075,124076,124077,124078,124079,124080,124081,124082,124083,124084,124085,124086,124087,124088,124089,124090,124091,124092,124093,124095,124096,124097,124098,124099,124100,124101,124102,124103,124104,124105,124106,124107,124108,124109,124110,124111,124112,124113,124114,124115,124116,124117,124118,124119,124120,124121,124122,124123,124124,124126,124127,124128,124129,124130,124131,124132,124133,124134,124135,124136,124137,124138,124139,124140,124141,124142,124143,124144,124145,124146,124147,124148,124149,124150,124151,124152,124153,124154,124155,124156,124157,124158,124159,124160,124161,124162,124163,124164,124165,124166,124167,124168,124169,124170,124171,124172,124173,124174,124175,124176,124177,124178,124179,124180,124181,124182,124183,124184,124185,124186,124186,124187,124188,124189,124190,124191,124192,124193,124194,124195,124196,124197,124198,124199,124200,124201,124202,124203,124204,124205,124206,124207,124208,124209,124210,124211,124212,124213,124214,124215,124216,124216,124217,124218,124219,124220,124221,124222,124223,124224,124225,124226,124227,124228,124229,124230,124231,124232,124233,124234,124235,124236,124236,124237,124238,124239,124240,124241,124242,124243,124244,124245,124246,124247,124248,124249,124250,124251,124251,124252,124253,124254,124255,124256,124257,124258,124259,124260,124261,124262,124263,124264,124264,124265,124266,124267,124268,124269,124270,124271,124272,124273,124274,124275,124276,124276,124277,124278,124279,124280,124281,124282,124283,124284,124285,124286,124286,124287,124288,124289,124290,124291,124292,124293,124294,124295,124296,124296,124297,124298,124299,124300,124301,124302,124303,124304,124305,124305,124306,124307,124308,124309,124310,124311,124312,124313,124314,124314,124315,124316,124317,124318,124319,124320,124321,124322,124322,124323,124324,124325,124326,124327,124328,124329,124329,124330,124331,124332,124333,124334,124335,124336,124337,124337,124338,124339,124340,124341,124342,124343,124344,124344,124345,124346,124347,124348,124349,124350,124350,124351,124352,124353,124354,124355,124356,124357,124357,124358,124359,124360,124361,124362,124363,124363,124364,124365,124366,124367,124368,124369,124369,124370,124371,124372,124373,124374,124375,124375,124376,124377,124378,124379,124380,124380,124381,124382,124383,124384,124385,124386,124386,124387,124388,124389,124390,124391,124391,124392,124393,124394,124395,124396,124397,124397,124398,124399,124400,124401,124402,124402,124403,124404,124405,124406,124407,124407,124408,124409,124410,124411,124412,124412,124413,124414,124415,124416,124416,124417,124418,124419,124420,124421,124421,124422,124423,124424,124425,124426,124426,124427,124428,124429,124430,124430,124431,124432,124433,124434,124434,124435,124436,124437,124438,124439,124439,124440,124441,124442,124443,124443,124444,124445,124446,124447,124447,124448,124449,124450,124451,124451,124452,124453,124454,124455,124455,124456,124457,124458,124459,124459,124460,124461,124462,124463,124463,124464,124465,124466,124467,124467,124468,124469,124470,124471,124471,124472,124473,124474,124475,124475,124476,124477,124478,124478,124479,124480,124481,124482,124482,124483,124484,124485,124486,124486,124487,124488,124489,124489,124490,124491,124492,124493,124493,124494,124495,124496,124496,124497,124498,124499,124500,124500,124501,124502,124503,124503,124504,124505,124506,124506,124507,124508,124509,124510,124510,124511,124512,124513,124513,124514,124515,124516,124516,124517,124518,124519,124519,124520,124521,124522,124522,124523,124524,124525,124526,124526,124527,124528,124529,124529,124530,124531,124532,124532,124533,124534,124535,124535,124536,124537,124538,124538,124539,124540,124541,124541,124542,124543,124544,124544,124545,124546,124547,124547,124548,124549,124549,124550,124551,124552,124552,124553,124554,124555,124555,124556,124557,124558,124558,124559,124560,124561,124561,124562,124563,124564,124564,124565,124566,124566,124567,124568,124569,124569,124570,124571,124572,124572,124573,124574,124574,124575,124576,124577,124577,124578,124579,124580,124580,124581,124582,124582,124583,124584,124585,124585,124586,124587,124587,124588,124589,124590,124590,124591,124592,124593,124593,124594,124595,124595,124596,124597,124598,124598,124599,124600,124600,124601,124602,124602,124603,124604,124605,124605,124606,124607,124607,124608,124609,124610,124610,124611,124612,124612,124613,124614,124615,124615,124616,124617,124617,124618,124619,124619,124620,124621,124622,124622,124623,124624,124624,124625,124626,124626,124627,124628,124628,124629,124630,124631,124631,124632,124633,124633,124634,124635,124635,124636,124637,124637,124638,124639,124640,124640,124641,124642,124642,124643,124644,124644,124645,124646,124646,124647,124648,124648,124649,124650,124651,124651,124652,124653,124653,124654,124655,124655,124656,124657,124657,124658,124659,124659,124660,124661,124661,124662,124663,124663,124664,124665,124665,124666,124667,124667,124668,124669,124669,124670,124671,124671,124672,124673,124674,124674,124675,124676,124676,124677,124678,124678,124679,124680,124680,124681,124682,124682,124683,124683,124684,124685,124685,124686,124687,124687,124688,124689,124689,124690,124691,124691,124692,124693,124693,124694,124695,124695,124696,124697,124697,124698,124699,124699,124700,124701,124701,124702,124703,124703,124704,124705,124705,124706,124706,124707,124708,124708,124709,124710,124710,124711,124712,124712,124713,124714,124714,124715,124716,124716,124717,124717,124718,124719,124719,124720,124721,124721,124722,124723,124723,124724,124725,124725,124726,124726,124727,124728,124728,124729,124730,124730,124731,124732,124732,124733,124733,124734,124735,124735,124736,124737,124737,124738,124739,124739,124740,124740,124741,124742,124742,124743,124744,124744,124745,124745,124746,124747,124747,124748,124749,124749,124750,124750,124751,124752,124752,124753,124754,124754,124755,124755,124756,124757,124757,124758,124759,124759,124760,124760,124761,124762,124762,124763,124764,124764,124765,124765,124766,124767,124767,124768,124768,124769,124770,124770,124771,124772,124772,124773,124773,124774,124775,124775,124776,124776,124777,124778,124778,124779,124779,124780,124781,124781,124782,124783,124783,124784,124784,124785,124786,124786,124787,124787,124788,124789,124789,124790,124790,124791,124792,124792,124793,124793,124794,124795,124795,124796,124796,124797,124798,124798,124799,124799,124800,124801,124801,124802,124802,124803,124804,124804,124805,124805,124806,124807,124807,124808,124808,124809,124810,124810,124811,124811,124812,124813,124813,124814,124814,124815,124815,124816,124817,124817,124818,124818,124819,124820,124820,124821,124821,124822,124823,124823,124824,124824,124825,124825,124826,124827,124827,124828,124828,124829,124830,124830,124831,124831,124832,124832,124833,124834,124834,124835,124835,124836,124836,124837,124838,124838,124839,124839,124840,124841,124841,124842,124842,124843,124843,124844,124845,124845,124846,124846,124847,124847,124848,124849,124849,124850,124850,124851,124851,124852,124853,124853,124854,124854,124855,124855,124856,124857,124857,124858,124858,124859,124859,124860,124861,124861,124862,124862,124863,124863,124864,124864,124865,124866,124866,124867,124867,124868,124868,124869,124870,124870,124871,124871,124872,124872,124873,124873,124874,124875,124875,124876,124876,124877,124877,124878,124878,124879,124880,124880,124881,124881,124882,124882,124883,124883,124884,124885,124885,124886,124886,124887,124887,124888,124888,124889,124890,124890,124891,124891,124892,124892,124893,124893,124894,124894,124895,124896,124896,124897,124897,124898,124898,124899,124899,124900,124900,124901,124902,124902,124903,124903,124904,124904,124905,124905,124906,124906,124907,124908,124908,124909,124909,124910,124910,124911,124911,124912,124912,124913,124913,124914,124915,124915,124916,124916,124917,124917,124918,124918,124919,124919,124920,124920,124921,124922,124922,124923,124923,124924,124924,124925,124925,124926,124926,124927,124927,124928,124928,124929,124930,124930,124931,124931,124932,124932,124933,124933,124934,124934,124935,124935,124936,124936,124937,124937,124938,124938,124939,124940,124940,124941,124941,124942,124942,124943,124943,124944,124944,124945,124945,124946,124946,124947,124947,124948,124948,124949,124949,124950,124950,124951,124952,124952,124953,124953,124954,124954,124955,124955,124956,124956,124957,124957,124958,124958,124959,124959,124960,124960,124961,124961,124962,124962,124963,124963,124964,124964,124965,124965,124966,124966,124967,124967,124968,124969,124969,124970,124970,124971,124971,124972,124972,124973,124973,124974,124974,124975,124975,124976,124976,124977,124977,124978,124978,124979,124979,124980,124980,124981,124981,124982,124982,124983,124983,124984,124984,124985,124985,124986,124986,124987,124987,124988,124988,124989,124989,124990,124990,124991,124991,124992,124992,124993,124993,124994,124994,124995,124995,124996,124996,124997,124997,124998,124998,124999,124999,125000,125000,125001,125001,125002,125002,125003,125003,125004,125004,125005,125005,125006,125006,125007,125007,125008,125008,125009,125009,125009,125010,125010,125011,125011,125012,125012,125013,125013,125014,125014,125015,125015,125016,125016,125017,125017,125018,125018,125019,125019,125020,125020,125021,125021,125022,125022,125023,125023,125024,125024,125025,125025,125026,125026,125026,125027,125027,125028,125028,125029,125029,125030,125030,125031,125031,125032,125032,125033,125033,125034,125034,125035,125035,125036,125036,125037,125037,125037,125038,125038,125039,125039,125040,125040,125041,125041,125042,125042,125043,125043,125044,125044,125045,125045,125046,125046,125046,125047,125047,125048,125048,125049,125049,125050,125050,125051,125051,125052,125052,125053,125053,125054,125054,125054,125055,125055,125056,125056,125057,125057,125058,125058,125059,125059,125060,125060,125061,125061,125061,125062,125062,125063,125063,125064,125064,125065,125065,125066,125066,125067,125067,125067,125068,125068,125069,125069,125070,125070,125071,125071,125072,125072,125073,125073,125073,125074,125074,125075,125075,125076,125076,125077,125077,125078,125078,125079,125079,125079,125080,125080,125081,125081,125082,125082,125083,125083,125084,125084,125084,125085,125085,125086,125086,125087,125087,125088,125088,125088,125089,125089,125090,125090,125091,125091,125092,125092,125093,125093,125093,125094,125094,125095,125095,125096,125096,125097,125097,125097,125098,125098,125099,125099,125100,125100,125101,125101,125101,125102,125102,125103,125103,125104,125104,125105,125105,125105,125106,125106,125107,125107,125108,125108,125109,125109,125109,125110,125110,125111,125111,125112,125112,125113,125113,125113,125114,125114,125115,125115,125116,125116,125117,125117,125117,125118,125118,125119,125119,125120,125120,125120,125121,125121,125122,125122,125123,125123,125124,125124,125124,125125,125125,125126,125126,125127,125127,125127,125128,125128,125129,125129,125130,125130,125130,125131,125131,125132,125132,125133,125133,125133,125134,125134,125135,125135,125136,125136,125136,125137,125137,125138,125138,125139,125139,125139,125140,125140,125141,125141,125142,125142,125142,125143,125143,125144,125144,125145,125145,125145,125146,125146,125147,125147,125148,125148,125148,125149,125149,125150,125150,125151,125151,125151,125152,125152,125153,125153,125153,125154,125154,125155,125155,125156,125156,125156,125157,125157,125158,125158,125159,125159,125159,125160,125160,125161,125161,125161,125162,125162,125163,125163,125164,125164,125164,125165,125165,125166,125166,125166,125167,125167,125168,125168,125169,125169,125169,125170,125170,125171,125171,125171,125172,125172,125173,125173,125174,125174,125174,125175,125175,125176,125176,125176,125177,125177,125178,125178,125178,125179,125179,125180,125180,125180,125181,125181,125182,125182,125183,125183,125183,125184,125184,125185,125185,125185,125186,125186,125187,125187,125187,125188,125188,125189,125189,125189,125190,125190,125191,125191,125191,125192,125192,125193,125193,125193,125194,125194,125195,125195,125195,125196,125196,125197,125197,125198,125198,125198,125199,125199,125200,125200,125200,125201,125201,125202,125202,125202,125203,125203,125204,125204,125204,125205,125205,125206,125206,125206,125207,125207,125207,125208,125208,125209,125209,125209,125210,125210,125211,125211,125211,125212,125212,125213,125213,125213,125214,125214,125215,125215,125215,125216,125216,125217,125217,125217,125218,125218,125219,125219,125219,125220,125220,125221,125221,125221,125222,125222,125222,125223,125223,125224,125224,125224,125225,125225,125226,125226,125226,125227,125227,125228,125228,125228,125229,125229,125229,125230,125230,125231,125231,125231,125232,125232,125233,125233,125233,125234,125234,125234,125235,125235,125236,125236,125236,125237,125237,125238,125238,125238,125239,125239,125239,125240,125240,125241,125241,125241,125242,125242,125243,125243,125243,125244,125244,125244,125245,125245,125246,125246,125246,125247,125247,125247,125248,125248,125249,125249,125249,125250,125250,125251,125251,125251,125252,125252,125252,125253,125253,125254,125254,125254,125255,125255,125255,125256,125256,125257,125257,125257,125258,125258,125258,125259,125259,125260,125260,125260,125261,125261,125261,125262,125262,125263,125263,125263,125264,125264,125264,125265,125265,125266,125266,125266,125267,125267,125267,125268,125268,125268,125269,125269,125270,125270,125270,125271,125271,125271,125272,125272,125273,125273,125273,125274,125274,125274,125275,125275,125275,125276,125276,125277,125277,125277,125278,125278,125278,125279,125279,125280,125280,125280,125281,125281,125281,125282,125282,125282,125283,125283,125284,125284,125284,125285,125285,125285,125286,125286,125286,125287,125287,125288,125288,125288,125289,125289,125289,125290,125290,125290,125291,125291,125292,125292,125292,125293,125293,125293,125294,125294,125294,125295,125295,125295,125296,125296,125297,125297,125297,125298,125298,125298,125299,125299,125299,125300,125300,125300,125301,125301,125302,125302,125302,125303,125303,125303,125304,125304,125304,125305,125305,125305,125306,125306,125307,125307,125307,125308,125308,125308,125309,125309,125309,125310,125310,125310,125311,125311,125311,125312,125312,125313,125313,125313,125314,125314,125314,125315,125315,125315,125316,125316,125316,125317,125317,125317,125318,125318,125319,125319,125319,125320,125320,125320,125321,125321,125321,125322,125322,125322,125323,125323,125323,125324,125324,125324,125325,125325,125325,125326,125326,125327,125327,125327,125328,125328,125328,125329,125329,125329,125330,125330,125330,125331,125331,125331,125332,125332,125332,125333,125333,125333,125334,125334,125334,125335,125335,125335,125336,125336,125336,125337,125337,125338,125338,125338,125339,125339,125339,125340,125340,125340,125341,125341,125341,125342,125342,125342,125343,125343,125343,125344,125344,125344,125345,125345,125345,125346,125346,125346,125347,125347,125347,125348,125348,125348,125349,125349,125349,125350,125350,125350,125351,125351,125351,125352,125352,125352,125353,125353,125353,125354,125354,125354,125355,125355,125355,125356,125356,125356,125357,125357,125357,125358,125358,125358,125359,125359,125359,125360,125360,125360,125361,125361,125361,125362,125362,125362,125363,125363,125363,125364,125364,125364,125365,125365,125365,125366,125366,125366,125367,125367,125367,125368,125368,125368,125369,125369,125369,125370,125370,125370,125371,125371,125371,125372,125372,125372,125373,125373,125373,125374,125374,125374,125375,125375,125375,125376,125376,125376,125377,125377,125377,125378,125378,125378,125378,125379,125379,125379,125380,125380,125380,125381,125381,125381,125382,125382,125382,125383,125383,125383,125384,125384,125384,125385,125385,125385,125386,125386,125386,125387,125387,125387,125388,125388,125388,125388,125389,125389,125389,125390,125390,125390,125391,125391,125391,125392,125392,125392,125393,125393,125393,125394,125394,125394,125395,125395,125395,125396,125396,125396,125396,125397,125397,125397,125398,125398,125398,125399,125399,125399,125400,125400,125400,125401,125401,125401,125402,125402,125402,125402,125403,125403,125403,125404,125404,125404,125405,125405,125405,125406,125406,125406,125407,125407,125407,125408,125408,125408,125408,125409,125409,125409,125410,125410,125410,125411,125411,125411,125412,125412,125412,125413,125413,125413,125413,125414,125414,125414,125415,125415,125415,125416,125416,125416,125417,125417,125417,125417,125418,125418,125418,125419,125419,125419,125420,125420,125420,125421,125421,125421,125422,125422,125422,125422,125423,125423,125423,125424,125424,125424,125425,125425,125425,125426,125426,125426,125426,125427,125427,125427,125428,125428,125428,125429,125429,125429,125429,125430,125430,125430,125431,125431,125431,125432,125432,125432,125433,125433,125433,125433,125434,125434,125434,125435,125435,125435,125436,125436,125436,125436,125437,125437,125437,125438,125438,125438,125439,125439,125439,125439,125440,125440,125440,125441,125441,125441,125442,125442,125442,125442,125443,125443,125443,125444,125444,125444,125445,125445,125445,125445,125446,125446,125446,125447,125447,125447,125448,125448,125448,125448,125449,125449,125449,125450,125450,125450,125451,125451,125451,125451,125452,125452,125452,125453,125453,125453,125453,125454,125454,125454,125455,125455,125455,125456,125456,125456,125456,125457,125457,125457,125458,125458,125458,125458,125459,125459,125459,125460,125460,125460,125461,125461,125461,125461,125462,125462,125462,125463,125463,125463,125463,125464,125464,125464,125465,125465,125465,125466,125466,125466,125466,125467,125467,125467,125468,125468,125468,125468,125469,125469,125469,125470,125470,125470,125470,125471,125471,125471,125472,125472,125472,125472,125473,125473,125473,125474,125474,125474,125474,125475,125475,125475,125476,125476,125476,125476,125477,125477,125477,125478,125478,125478,125478,125479,125479,125479,125480,125480,125480,125480,125481,125481,125481,125482,125482,125482,125482,125483,125483,125483,125484,125484,125484,125484,125485,125485,125485,125486,125486,125486,125486,125487,125487,125487,125488,125488,125488,125488,125489,125489,125489,125490,125490,125490,125490,125491,125491,125491,125492,125492,125492,125492,125493,125493,125493,125494,125494,125494,125494,125495,125495,125495,125495,125496,125496,125496,125497,125497,125497,125497,125498,125498,125498,125499,125499,125499,125499,125500,125500,125500,125500,125501,125501,125501,125502,125502,125502,125502,125503,125503,125503,125504,125504,125504,125504,125505,125505,125505,125505,125506,125506,125506,125507,125507,125507,125507,125508,125508,125508,125509,125509,125509,125509,125510,125510,125510,125510,125511,125511,125511,125512,125512,125512,125512,125513,125513,125513,125513,125514,125514,125514,125515,125515,125515,125515,125516,125516,125516,125516,125517,125517,125517,125518,125518,125518,125518,125519,125519,125519,125519,125520,125520,125520,125521,125521,125521,125521,125522,125522,125522,125522,125523,125523,125523,125523,125524,125524,125524,125525,125525,125525,125525,125526,125526,125526,125526,125527,125527,125527,125528,125528,125528,125528,125529,125529,125529,125529,125530,125530,125530,125530,125531,125531,125531,125532,125532,125532,125532,125533,125533,125533,125533,125534,125534,125534,125534,125535,125535,125535,125536,125536,125536,125536,125537,125537,125537,125537,125538,125538,125538,125538,125539,125539,125539,125539,125540,125540,125540,125541,125541,125541,125541,125542,125542,125542,125542,125543,125543,125543,125543,125544,125544,125544,125544,125545,125545,125545,125546,125546,125546,125546,125547,125547,125547,125547,125548,125548,125548,125548,125549,125549,125549,125549,125550,125550,125550,125550,125551,125551,125551,125551,125552,125552,125552,125553,125553,125553,125553,125554,125554,125554,125554,125555,125555,125555,125555,125556,125556,125556,125556,125557,125557,125557,125557,125558,125558,125558,125558,125559,125559,125559,125559,125560,125560,125560,125561,125561,125561,125561,125562,125562,125562,125562,125563,125563,125563,125563,125564,125564,125564,125564,125565,125565,125565,125565,125566,125566,125566,125566,125567,125567,125567,125567,125568,125568,125568,125568,125569,125569,125569,125569,125570,125570,125570,125570,125571,125571,125571,125571,125572,125572,125572,125572,125573,125573,125573,125573,125574,125574,125574,125574,125575,125575,125575,125575,125576,125576,125576,125576,125577,125577,125577,125577,125578,125578,125578,125578,125579,125579,125579,125579,125580,125580,125580,125580,125581,125581,125581,125581,125582,125582,125582,125582,125583,125583,125583,125583,125584,125584,125584,125584,125585,125585,125585,125585,125586,125586,125586,125586,125587,125587,125587,125587,125588,125588,125588,125588,125589,125589,125589,125589,125590,125590,125590,125590,125591,125591,125591,125591,125592,125592,125592,125592,125593,125593,125593,125593,125594,125594,125594,125594,125595,125595,125595,125595,125595,125596,125596,125596,125596,125597,125597,125597,125597,125598,125598,125598,125598,125599,125599,125599,125599,125600,125600,125600,125600,125601,125601,125601,125601,125602,125602,125602,125602,125603,125603,125603,125603,125603,125604,125604,125604,125604,125605,125605,125605,125605,125606,125606,125606,125606,125607,125607,125607,125607,125608,125608,125608,125608,125609,125609,125609,125609,125609,125610,125610,125610,125610,125611,125611,125611,125611,125612,125612,125612,125612,125613,125613,125613,125613,125614,125614,125614,125614,125614,125615,125615,125615,125615,125616,125616,125616,125616,125617,125617,125617,125617,125618,125618,125618,125618,125619,125619,125619,125619,125619,125620,125620,125620,125620,125621,125621,125621,125621,125622,125622,125622,125622,125623,125623,125623,125623,125623,125624,125624,125624,125624,125625,125625,125625,125625,125626,125626,125626,125626,125626,125627,125627,125627,125627,125628,125628,125628,125628,125629,125629,125629,125629,125630,125630,125630,125630,125630,125631,125631,125631,125631,125632,125632,125632,125632,125633,125633,125633,125633,125633,125634,125634,125634,125634,125635,125635,125635,125635,125636,125636,125636,125636,125636,125637,125637,125637,125637,125638,125638,125638,125638,125639,125639,125639,125639,125639,125640,125640,125640,125640,125641,125641,125641,125641,125641,125642,125642,125642,125642,125643,125643,125643,125643,125644,125644,125644,125644,125644,125645,125645,125645,125645,125646,125646,125646,125646,125646,125647,125647,125647,125647,125648,125648,125648,125648,125649,125649,125649,125649,125649,125650,125650,125650,125650,125651,125651,125651,125651,125651,125652,125652,125652,125652,125653,125653,125653,125653,125653,125654,125654,125654,125654,125655,125655,125655,125655,125655,125656,125656,125656,125656,125657,125657,125657,125657,125657,125658,125658,125658,125658,125659,125659,125659,125659,125659,125660,125660,125660,125660,125661,125661,125661,125661,125661,125662,125662,125662,125662,125663,125663,125663,125663,125663,125664,125664,125664,125664,125665,125665,125665,125665,125665,125666,125666,125666,125666,125667,125667,125667,125667,125667,125668,125668,125668,125668,125669,125669,125669,125669,125669,125670,125670,125670,125670,125670,125671,125671,125671,125671,125672,125672,125672,125672,125672,125673,125673,125673,125673,125674,125674,125674,125674,125674,125675,125675,125675,125675,125675,125676,125676,125676,125676,125677,125677,125677,125677,125677,125678,125678,125678,125678,125679,125679,125679,125679,125679,125680,125680,125680,125680,125680,125681,125681,125681,125681,125682,125682,125682,125682,125682,125683,125683,125683,125683,125683,125684,125684,125684,125684,125685,125685,125685,125685,125685,125686,125686,125686,125686,125686,125687,125687,125687,125687,125688,125688,125688,125688,125688,125689,125689,125689,125689,125689,125690,125690,125690,125690,125691,125691,125691,125691,125691,125692,125692,125692,125692,125692,125693,125693,125693,125693,125693,125694,125694,125694,125694,125695,125695,125695,125695,125695,125696,125696,125696,125696,125696,125697,125697,125697,125697,125697,125698,125698,125698,125698,125699,125699,125699,125699,125699,125700,125700,125700,125700,125700,125701,125701,125701,125701,125701,125702,125702,125702,125702,125702,125703,125703,125703,125703,125704,125704,125704,125704,125704,125705,125705,125705,125705,125705,125706,125706,125706,125706,125706,125707,125707,125707,125707,125707,125708,125708,125708,125708,125708,125709,125709,125709,125709,125710,125710,125710,125710,125710,125711,125711,125711,125711,125711,125712,125712,125712,125712,125712,125713,125713,125713,125713,125713,125714,125714,125714,125714,125714,125715,125715,125715,125715,125715,125716,125716,125716,125716,125716,125717,125717,125717,125717,125717,125718,125718,125718,125718,125718,125719,125719,125719,125719,125720,125720,125720,125720,125720,125721,125721,125721,125721,125721,125722,125722,125722,125722,125722,125723,125723,125723,125723,125723,125724,125724,125724,125724,125724,125725,125725,125725,125725,125725,125726,125726,125726,125726,125726,125727,125727,125727,125727,125727,125728,125728,125728,125728,125728,125729,125729,125729,125729,125729,125730,125730,125730,125730,125730,125731,125731,125731,125731,125731,125732,125732,125732,125732,125732,125733,125733,125733,125733,125733,125734,125734,125734,125734,125734,125735,125735,125735,125735,125735,125736,125736,125736,125736,125736,125737,125737,125737,125737,125737,125737,125738,125738,125738,125738,125738,125739,125739,125739,125739,125739,125740,125740,125740,125740,125740,125741,125741,125741,125741,125741,125742,125742,125742,125742,125742,125743,125743,125743,125743,125743,125744,125744,125744,125744,125744,125745,125745,125745,125745,125745,125746,125746,125746,125746,125746,125746,125747,125747,125747,125747,125747,125748,125748,125748,125748,125748,125749,125749,125749,125749,125749,125750,125750,125750,125750,125750,125751,125751,125751,125751,125751,125752,125752,125752,125752,125752,125752,125753,125753,125753,125753,125753,125754,125754,125754,125754,125754,125755,125755,125755,125755,125755,125756,125756,125756,125756,125756,125757,125757,125757,125757,125757,125757,125758,125758,125758,125758,125758,125759,125759,125759,125759,125759,125760,125760,125760,125760,125760,125761,125761,125761,125761,125761,125761,125762,125762,125762,125762,125762,125763,125763,125763,125763,125763,125764,125764,125764,125764,125764,125764,125765,125765,125765,125765,125765,125766,125766,125766,125766,125766,125767,125767,125767,125767,125767,125767,125768,125768,125768,125768,125768,125769,125769,125769,125769,125769,125770,125770,125770,125770,125770,125770,125771,125771,125771,125771,125771,125772,125772,125772,125772,125772,125773,125773,125773,125773,125773,125773,125774,125774,125774,125774,125774,125775,125775,125775,125775,125775,125776,125776,125776,125776,125776,125776,125777,125777,125777,125777,125777,125778,125778,125778,125778,125778,125778,125779,125779,125779,125779,125779,125780,125780,125780,125780,125780,125780,125781,125781,125781,125781,125781,125782,125782,125782,125782,125782,125783,125783,125783,125783,125783,125783,125784,125784,125784,125784,125784,125785,125785,125785,125785,125785,125785,125786,125786,125786,125786,125786,125787,125787,125787,125787,125787,125787,125788,125788,125788,125788,125788,125789,125789,125789,125789,125789,125789,125790,125790,125790,125790,125790,125791,125791,125791,125791,125791,125791,125792,125792,125792,125792,125792,125793,125793,125793,125793,125793,125793,125794,125794,125794,125794,125794,125794,125795,125795,125795,125795,125795,125796,125796,125796,125796,125796,125796,125797,125797,125797,125797,125797,125798,125798,125798,125798,125798,125798,125799,125799,125799,125799,125799,125799,125800,125800,125800,125800,125800,125801,125801,125801,125801,125801,125801,125802,125802,125802,125802,125802,125803,125803,125803,125803,125803,125803,125804,125804,125804,125804,125804,125804,125805,125805,125805,125805,125805,125806,125806,125806,125806,125806,125806,125807,125807,125807,125807,125807,125807,125808,125808,125808,125808,125808,125809,125809,125809,125809,125809,125809,125810,125810,125810,125810,125810,125810,125811,125811,125811,125811,125811,125811,125812,125812,125812,125812,125812,125813,125813,125813,125813,125813,125813,125814,125814,125814,125814,125814,125814,125815,125815,125815,125815,125815,125815,125816,125816,125816,125816,125816,125817,125817,125817,125817,125817,125817,125818,125818,125818,125818,125818,125818,125819,125819,125819,125819,125819,125819,125820,125820,125820,125820,125820,125820,125821,125821,125821,125821,125821,125822,125822,125822,125822,125822,125822,125823,125823,125823,125823,125823,125823,125824,125824,125824,125824,125824,125824,125825,125825,125825,125825,125825,125825,125826,125826,125826,125826,125826,125826,125827,125827,125827,125827,125827,125827,125828,125828,125828,125828,125828,125829,125829,125829,125829,125829,125829,125830,125830,125830,125830,125830,125830,125831,125831,125831,125831,125831,125831,125832,125832,125832,125832,125832,125832,125833,125833,125833,125833,125833,125833,125834,125834,125834,125834,125834,125834,125835,125835,125835,125835,125835,125835,125836,125836,125836,125836,125836,125836,125837,125837,125837,125837,125837,125837,125838,125838,125838,125838,125838,125838,125839,125839,125839,125839,125839,125839,125840,125840,125840,125840,125840,125840,125841,125841,125841,125841,125841,125841,125842,125842,125842,125842,125842,125842,125843,125843,125843,125843,125843,125843,125844,125844,125844,125844,125844,125844,125845,125845,125845,125845,125845,125845,125846,125846,125846,125846,125846,125846,125847,125847,125847,125847,125847,125847,125848,125848,125848,125848,125848,125848,125849,125849,125849,125849,125849,125849,125849,125850,125850,125850,125850,125850,125850,125851,125851,125851,125851,125851,125851,125852,125852,125852,125852,125852,125852,125853,125853,125853,125853,125853,125853,125854,125854,125854,125854,125854,125854,125855,125855,125855,125855,125855,125855,125856,125856,125856,125856,125856,125856,125856,125857,125857,125857,125857,125857,125857,125858,125858,125858,125858,125858,125858,125859,125859,125859,125859,125859,125859,125860,125860,125860,125860,125860,125860,125861,125861,125861,125861,125861,125861,125861,125862,125862,125862,125862,125862,125862,125863,125863,125863,125863,125863,125863,125864,125864,125864,125864,125864,125864,125865,125865,125865,125865,125865,125865,125865,125866,125866,125866,125866,125866,125866,125867,125867,125867,125867,125867,125867,125868,125868,125868,125868,125868,125868,125868,125869,125869,125869,125869,125869,125869,125870,125870,125870,125870,125870,125870,125871,125871,125871,125871,125871,125871,125871,125872,125872,125872,125872,125872,125872,125873,125873,125873,125873,125873,125873,125874,125874,125874,125874,125874,125874,125874,125875,125875,125875,125875,125875,125875,125876,125876,125876,125876,125876,125876,125876,125877,125877,125877,125877,125877,125877,125878,125878,125878,125878,125878,125878,125879,125879,125879,125879,125879,125879,125879,125880,125880,125880,125880,125880,125880,125881,125881,125881,125881,125881,125881,125881,125882,125882,125882,125882,125882,125882,125883,125883,125883,125883,125883,125883,125883,125884,125884,125884,125884,125884,125884,125885,125885,125885,125885,125885,125885,125885,125886,125886,125886,125886,125886,125886,125887,125887,125887,125887,125887,125887,125887,125888,125888,125888,125888,125888,125888,125889,125889,125889,125889,125889,125889,125889,125890,125890,125890,125890,125890,125890,125891,125891,125891,125891,125891,125891,125891,125892,125892,125892,125892,125892,125892,125892,125893,125893,125893,125893,125893,125893,125894,125894,125894,125894,125894,125894,125894,125895,125895,125895,125895,125895,125895,125896,125896,125896,125896,125896,125896,125896,125897,125897,125897,125897,125897,125897,125897,125898,125898,125898,125898,125898,125898,125899,125899,125899,125899,125899,125899,125899,125900,125900,125900,125900,125900,125900,125900,125901,125901,125901,125901,125901,125901,125901,125902,125902,125902,125902,125902,125902,125903,125903,125903,125903,125903,125903,125903,125904,125904,125904,125904,125904,125904,125904,125905,125905,125905,125905,125905,125905,125906,125906,125906,125906,125906,125906,125906,125907,125907,125907,125907,125907,125907,125907,125908,125908,125908,125908,125908,125908,125908,125909,125909,125909,125909,125909,125909,125909,125910,125910,125910,125910,125910,125910,125911,125911,125911,125911,125911,125911,125911,125912,125912,125912,125912,125912,125912,125912,125913,125913,125913,125913,125913,125913,125913,125914,125914,125914,125914,125914,125914,125914,125915,125915,125915,125915,125915,125915,125915,125916,125916,125916,125916,125916,125916,125917,125917,125917,125917,125917,125917,125917,125918,125918,125918,125918,125918,125918,125918,125919,125919,125919,125919,125919,125919,125919,125920,125920,125920,125920,125920,125920,125920,125921,125921,125921,125921,125921,125921,125921,125922,125922,125922,125922,125922,125922,125922,125923,125923,125923,125923,125923,125923,125923,125924,125924,125924,125924,125924,125924,125924,125925,125925,125925,125925,125925,125925,125925,125926,125926,125926,125926,125926,125926,125926,125927,125927,125927,125927,125927,125927,125927,125928,125928,125928,125928,125928,125928,125928,125929,125929,125929,125929,125929,125929,125929,125930,125930,125930,125930,125930,125930,125930,125931,125931,125931,125931,125931,125931,125931,125932,125932,125932,125932,125932,125932,125932,125933,125933,125933,125933,125933,125933,125933,125933,125934,125934,125934,125934,125934,125934,125934,125935,125935,125935,125935,125935,125935,125935,125936,125936,125936,125936,125936,125936,125936,125937,125937,125937,125937,125937,125937,125937,125938,125938,125938,125938,125938,125938,125938,125939,125939,125939,125939,125939,125939,125939,125940,125940,125940,125940,125940,125940,125940,125940,125941,125941,125941,125941,125941,125941,125941,125942,125942,125942,125942,125942,125942,125942,125943,125943,125943,125943,125943,125943,125943,125944,125944,125944,125944,125944,125944,125944,125944,125945,125945,125945,125945,125945,125945,125945,125946,125946,125946,125946,125946,125946,125946,125947,125947,125947,125947,125947,125947,125947,125948,125948,125948,125948,125948,125948,125948,125948,125949,125949,125949,125949,125949,125949,125949,125950,125950,125950,125950,125950,125950,125950,125951,125951,125951,125951,125951,125951,125951,125951,125952,125952,125952,125952,125952,125952,125952,125953,125953,125953,125953,125953,125953,125953,125953,125954,125954,125954,125954,125954,125954,125954,125955,125955,125955,125955,125955,125955,125955,125956,125956,125956,125956,125956,125956,125956,125956,125957,125957,125957,125957,125957,125957,125957,125958,125958,125958,125958,125958,125958,125958,125958,125959,125959,125959,125959,125959,125959,125959,125960,125960,125960,125960,125960,125960,125960,125960,125961,125961,125961,125961,125961,125961,125961,125962,125962,125962,125962,125962,125962,125962,125962,125963,125963,125963,125963,125963,125963,125963,125964,125964,125964,125964,125964,125964,125964,125964,125965,125965,125965,125965,125965,125965,125965,125966,125966,125966,125966,125966,125966,125966,125966,125967,125967,125967,125967,125967,125967,125967,125968,125968,125968,125968,125968,125968,125968,125968,125969,125969,125969,125969,125969,125969,125969,125969,125970,125970,125970,125970,125970,125970,125970,125971,125971,125971,125971,125971,125971,125971,125971,125972,125972,125972,125972,125972,125972,125972,125972,125973,125973,125973,125973,125973,125973,125973,125974,125974,125974,125974,125974,125974,125974,125974,125975,125975,125975,125975,125975,125975,125975,125975,125976,125976,125976,125976,125976,125976,125976,125977,125977,125977,125977,125977,125977,125977,125977,125978,125978,125978,125978,125978,125978,125978,125978,125979,125979,125979,125979,125979,125979,125979,125979,125980,125980,125980,125980,125980,125980,125980,125981,125981,125981,125981,125981,125981,125981,125981,125982,125982,125982,125982,125982,125982,125982,125982,125983,125983,125983,125983,125983,125983,125983,125983,125984,125984,125984,125984,125984,125984,125984,125984,125985,125985,125985,125985,125985,125985,125985,125985,125986,125986,125986,125986,125986,125986,125986,125987,125987,125987,125987,125987,125987,125987,125987,125988,125988,125988,125988,125988,125988,125988,125988,125989,125989,125989,125989,125989,125989,125989,125989,125990,125990,125990,125990,125990,125990,125990,125990,125991,125991,125991,125991,125991,125991,125991,125991,125992,125992,125992,125992,125992,125992,125992,125992,125993,125993,125993,125993,125993,125993,125993,125993,125994,125994,125994,125994,125994,125994,125994,125994,125995,125995,125995,125995,125995,125995,125995,125995,125996,125996,125996,125996,125996,125996,125996,125996,125997,125997,125997,125997,125997,125997,125997,125997,125998,125998,125998,125998,125998,125998,125998,125998,125999,125999,125999,125999,125999,125999,125999,125999,126000,126000,126000,126000,126000,126000,126000,126000,126001,126001,126001,126001,126001,126001,126001,126001,126002,126002,126002,126002,126002,126002,126002,126002,126003,126003,126003,126003,126003,126003,126003,126003,126003,126004,126004,126004,126004,126004,126004,126004,126004,126005,126005,126005,126005,126005,126005,126005,126005,126006,126006,126006,126006,126006,126006,126006,126006,126007,126007,126007,126007,126007,126007,126007,126007,126008,126008,126008,126008,126008,126008,126008,126008,126008,126009,126009,126009,126009,126009,126009,126009,126009,126010,126010,126010,126010,126010,126010,126010,126010,126011,126011,126011,126011,126011,126011,126011,126011,126012,126012,126012,126012,126012,126012,126012,126012,126012,126013,126013,126013,126013,126013,126013,126013,126013,126014,126014,126014,126014,126014,126014,126014,126014,126015,126015,126015,126015,126015,126015,126015,126015,126015,126016,126016,126016,126016,126016,126016,126016,126016,126017,126017,126017,126017,126017,126017,126017,126017,126018,126018,126018,126018,126018,126018,126018,126018,126018,126019,126019,126019,126019,126019,126019,126019,126019,126020,126020,126020,126020,126020,126020,126020,126020,126020,126021,126021,126021,126021,126021,126021,126021,126021,126022,126022,126022,126022,126022,126022,126022,126022,126022,126023,126023,126023,126023,126023,126023,126023,126023,126024,126024,126024,126024,126024,126024,126024,126024,126025,126025,126025,126025,126025,126025,126025,126025,126025,126026,126026,126026,126026,126026,126026,126026,126026,126026,126027,126027,126027,126027,126027,126027,126027,126027,126028,126028,126028,126028,126028,126028,126028,126028,126028,126029,126029,126029,126029,126029,126029,126029,126029,126030,126030,126030,126030,126030,126030,126030,126030,126030,126031,126031,126031,126031,126031,126031,126031,126031,126032,126032,126032,126032,126032,126032,126032,126032,126032,126033,126033,126033,126033,126033,126033,126033,126033,126033,126034,126034,126034,126034,126034,126034,126034,126034,126035,126035,126035,126035,126035,126035,126035,126035,126035,126036,126036,126036,126036,126036,126036,126036,126036,126036,126037,126037,126037,126037,126037,126037,126037,126037,126037,126038,126038,126038,126038,126038,126038,126038,126038,126039,126039,126039,126039,126039,126039,126039,126039,126039,126040,126040,126040,126040,126040,126040,126040,126040,126040,126041,126041,126041,126041,126041,126041,126041,126041,126041,126042,126042,126042,126042,126042,126042,126042,126042,126043,126043,126043,126043,126043,126043,126043,126043,126043,126044,126044,126044,126044,126044,126044,126044,126044,126044,126045,126045,126045,126045,126045,126045,126045,126045,126045,126046,126046,126046,126046,126046,126046,126046,126046,126046,126047,126047,126047,126047,126047,126047,126047,126047,126047,126048,126048,126048,126048,126048,126048,126048,126048,126048,126049,126049,126049,126049,126049,126049,126049,126049,126049,126050,126050,126050,126050,126050,126050,126050,126050,126050,126051,126051,126051,126051,126051,126051,126051,126051,126051,126052,126052,126052,126052,126052,126052,126052,126052,126052,126053,126053,126053,126053,126053,126053,126053,126053,126053,126054,126054,126054,126054,126054,126054,126054,126054,126054,126055,126055,126055,126055,126055,126055,126055,126055,126055,126056,126056,126056,126056,126056,126056,126056,126056,126056,126057,126057,126057,126057,126057,126057,126057,126057,126057,126058,126058,126058,126058,126058,126058,126058,126058,126058,126059,126059,126059,126059,126059,126059,126059,126059,126059,126060,126060,126060,126060,126060,126060,126060,126060,126060,126061,126061,126061,126061,126061,126061,126061,126061,126061,126061,126062,126062,126062,126062,126062,126062,126062,126062,126062,126063,126063,126063,126063,126063,126063,126063,126063,126063,126064,126064,126064,126064,126064,126064,126064,126064,126064,126065,126065,126065,126065,126065,126065,126065,126065,126065,126065,126066,126066,126066,126066,126066,126066,126066,126066,126066,126067,126067,126067,126067,126067,126067,126067,126067,126067,126068,126068,126068,126068,126068,126068,126068,126068,126068,126069,126069,126069,126069,126069,126069,126069,126069,126069,126069,126070,126070,126070,126070,126070,126070,126070,126070,126070,126071,126071,126071,126071,126071,126071,126071,126071,126071,126072,126072,126072,126072,126072,126072,126072,126072,126072,126072,126073,126073,126073,126073,126073,126073,126073,126073,126073,126074,126074,126074,126074,126074,126074,126074,126074,126074,126074,126075,126075,126075,126075,126075,126075,126075,126075,126075,126076,126076,126076,126076,126076,126076,126076,126076,126076,126076,126077,126077,126077,126077,126077,126077,126077,126077,126077,126078,126078,126078,126078,126078,126078,126078,126078,126078,126078,126079,126079,126079,126079,126079,126079,126079,126079,126079,126080,126080,126080,126080,126080,126080,126080,126080,126080,126080,126081,126081,126081,126081,126081,126081,126081,126081,126081,126082,126082,126082,126082,126082,126082,126082,126082,126082,126082,126083,126083,126083,126083,126083,126083,126083,126083,126083,126083,126084,126084,126084,126084,126084,126084,126084,126084,126084,126085,126085,126085,126085,126085,126085,126085,126085,126085,126085,126086,126086,126086,126086,126086,126086,126086,126086,126086,126086,126087,126087,126087,126087,126087,126087,126087,126087,126087,126088,126088,126088,126088,126088,126088,126088,126088,126088,126088,126089,126089,126089,126089,126089,126089,126089,126089,126089,126089,126090,126090,126090,126090,126090,126090,126090,126090,126090,126090,126091,126091,126091,126091,126091,126091,126091,126091,126091,126092,126092,126092,126092,126092,126092,126092,126092,126092,126092,126093,126093,126093,126093,126093,126093,126093,126093,126093,126093,126094,126094,126094,126094,126094,126094,126094,126094,126094,126094,126095,126095,126095,126095,126095,126095,126095,126095,126095,126095,126096,126096,126096,126096,126096,126096,126096,126096,126096,126096,126097,126097,126097,126097,126097,126097,126097,126097,126097,126097,126098,126098,126098,126098,126098,126098,126098,126098,126098,126098,126099,126099,126099,126099,126099,126099,126099,126099,126099,126099,126100,126100,126100,126100,126100,126100,126100,126100,126100,126100,126101,126101,126101,126101,126101,126101,126101,126101,126101,126101,126102,126102,126102,126102,126102,126102,126102,126102,126102,126102,126103,126103,126103,126103,126103,126103,126103,126103,126103,126103,126104,126104,126104,126104,126104,126104,126104,126104,126104,126104,126105,126105,126105,126105,126105,126105,126105,126105,126105,126105,126106,126106,126106,126106,126106,126106,126106,126106,126106,126106,126107,126107,126107,126107,126107,126107,126107,126107,126107,126107,126108,126108,126108,126108,126108,126108,126108,126108,126108,126108,126109,126109,126109,126109,126109,126109,126109,126109,126109,126109,126110,126110,126110,126110,126110,126110,126110,126110,126110,126110,126110,126111,126111,126111,126111,126111,126111,126111,126111,126111,126111,126112,126112,126112,126112,126112,126112,126112,126112,126112,126112,126113,126113,126113,126113,126113,126113,126113,126113,126113,126113,126114,126114,126114,126114,126114,126114,126114,126114,126114,126114,126114,126115,126115,126115,126115,126115,126115,126115,126115,126115,126115,126116,126116,126116,126116,126116,126116,126116,126116,126116,126116,126116,126117,126117,126117,126117,126117,126117,126117,126117,126117,126117,126118,126118,126118,126118,126118,126118,126118,126118,126118,126118,126119,126119,126119,126119,126119,126119,126119,126119,126119,126119,126119,126120,126120,126120,126120,126120,126120,126120,126120,126120,126120,126121,126121,126121,126121,126121,126121,126121,126121,126121,126121,126121,126122,126122,126122,126122,126122,126122,126122,126122,126122,126122,126123,126123,126123,126123,126123,126123,126123,126123,126123,126123,126123,126124,126124,126124,126124,126124,126124,126124,126124,126124,126124,126125,126125,126125,126125,126125,126125,126125,126125,126125,126125,126125,126126,126126,126126,126126,126126,126126,126126,126126,126126,126126,126127,126127,126127,126127,126127,126127,126127,126127,126127,126127,126127,126128,126128,126128,126128,126128,126128,126128,126128,126128,126128,126128,126129,126129,126129,126129,126129,126129,126129,126129,126129,126129,126130,126130,126130,126130,126130,126130,126130,126130,126130,126130,126130,126131,126131,126131,126131,126131,126131,126131,126131,126131,126131,126131,126132,126132,126132,126132,126132,126132,126132,126132,126132,126132,126133,126133,126133,126133,126133,126133,126133,126133,126133,126133,126133,126134,126134,126134,126134,126134,126134,126134,126134,126134,126134,126134,126135,126135,126135,126135,126135,126135,126135,126135,126135,126135,126135,126136,126136,126136,126136,126136,126136,126136,126136,126136,126136,126136,126137,126137,126137,126137,126137,126137,126137,126137,126137,126137,126137,126138,126138,126138,126138,126138,126138,126138,126138,126138,126138,126139,126139,126139,126139,126139,126139,126139,126139,126139,126139,126139,126140,126140,126140,126140,126140,126140,126140,126140,126140,126140,126140,126141,126141,126141,126141,126141,126141,126141,126141,126141,126141,126141,126142,126142,126142,126142,126142,126142,126142,126142,126142,126142,126142,126143,126143,126143,126143,126143,126143,126143,126143,126143,126143,126143,126144,126144,126144,126144,126144,126144,126144,126144,126144,126144,126144,126145,126145,126145,126145,126145,126145,126145,126145,126145,126145,126145,126146,126146,126146,126146,126146,126146,126146,126146,126146,126146,126146,126146,126147,126147,126147,126147,126147,126147,126147,126147,126147,126147,126147,126148,126148,126148,126148,126148,126148,126148,126148,126148,126148,126148,126149,126149,126149,126149,126149,126149,126149,126149,126149,126149,126149,126150,126150,126150,126150,126150,126150,126150,126150,126150,126150,126150,126151,126151,126151,126151,126151,126151,126151,126151,126151,126151,126151,126152,126152,126152,126152,126152,126152,126152,126152,126152,126152,126152,126152,126153,126153,126153,126153,126153,126153,126153,126153,126153,126153,126153,126154,126154,126154,126154,126154,126154,126154,126154,126154,126154,126154,126155,126155,126155,126155,126155,126155,126155,126155,126155,126155,126155,126155,126156,126156,126156,126156,126156,126156,126156,126156,126156,126156,126156,126157,126157,126157,126157,126157,126157,126157,126157,126157,126157,126157,126158,126158,126158,126158,126158,126158,126158,126158,126158,126158,126158,126158,126159,126159,126159,126159,126159,126159,126159,126159,126159,126159,126159,126160,126160,126160,126160,126160,126160,126160,126160,126160,126160,126160,126160,126161,126161,126161,126161,126161,126161,126161,126161,126161,126161,126161,126162,126162,126162,126162,126162,126162,126162,126162,126162,126162,126162,126162,126163,126163,126163,126163,126163,126163,126163,126163,126163,126163,126163,126164,126164,126164,126164,126164,126164,126164,126164,126164,126164,126164,126164,126165,126165,126165,126165,126165,126165,126165,126165,126165,126165,126165,126166,126166,126166,126166,126166,126166,126166,126166,126166,126166,126166,126166,126167,126167,126167,126167,126167,126167,126167,126167,126167,126167,126167,126167,126168,126168,126168,126168,126168,126168,126168,126168,126168,126168,126168,126169,126169,126169,126169,126169,126169,126169,126169,126169,126169,126169,126169,126170,126170,126170,126170,126170,126170,126170,126170,126170,126170,126170,126170,126171,126171,126171,126171,126171,126171,126171,126171,126171,126171,126171,126171,126172,126172,126172,126172,126172,126172,126172,126172,126172,126172,126172,126172,126173,126173,126173,126173,126173,126173,126173,126173,126173,126173,126173,126174,126174,126174,126174,126174,126174,126174,126174,126174,126174,126174,126174,126175,126175,126175,126175,126175,126175,126175,126175,126175,126175,126175,126175,126176,126176,126176,126176,126176,126176,126176,126176,126176,126176,126176,126176,126177,126177,126177,126177,126177,126177,126177,126177,126177,126177,126177,126177,126178,126178,126178,126178,126178,126178,126178,126178,126178,126178,126178,126178,126179,126179,126179,126179,126179,126179,126179,126179,126179,126179,126179,126179,126180,126180,126180,126180,126180,126180,126180,126180,126180,126180,126180,126180,126181,126181,126181,126181,126181,126181,126181,126181,126181,126181,126181,126181,126182,126182,126182,126182,126182,126182,126182,126182,126182,126182,126182,126182,126183,126183,126183,126183,126183,126183,126183,126183,126183,126183,126183,126183,126184,126184,126184,126184,126184,126184,126184,126184,126184,126184,126184,126184,126185,126185,126185,126185,126185,126185,126185,126185,126185,126185,126185,126185,126185,126186,126186,126186,126186,126186,126186,126186,126186,126186,126186,126186,126186,126187,126187,126187,126187,126187,126187,126187,126187,126187,126187,126187,126187,126188,126188,126188,126188,126188,126188,126188,126188,126188,126188,126188,126188,126189,126189,126189,126189,126189,126189,126189,126189,126189,126189,126189,126189,126189,126190,126190,126190,126190,126190,126190,126190,126190,126190,126190,126190,126190,126191,126191,126191,126191,126191,126191,126191);
        variable x       : integer := valores'length;
        variable valor   : integer := 127000;
    begin
        if ( z_accel /= 0 ) then
            x := abs(y_accel) * 100 / abs(z_accel);
        end if;
        if ( x < valores'length ) then
            valor := valores(x);
        end if;
        if y_accel < 0 then
            valor := -valor;
        end if;
        return valor;
    end calc_angulo_crudo;
        
begin

    process(reloj)
        variable x_gyro_integer      : integer;
        variable y_gyro_integer      : integer;
        variable y_accel_integer     : integer;
        variable z_accel_integer     : integer;
        variable angulo_crudo        : integer;
        variable omega_dt            : integer;
        variable angulo_filtrado     : integer := 0;
        variable velocidad           : integer;
        variable velocidad_fin       : integer;
        variable velocidad_a_temp    : integer;
        variable velocidad_b_temp    : integer;
        variable contador            : integer := 0;
        variable error               : integer := 0;
        variable dErr                : integer := 0;
        variable sum_error           : integer := 0;
        variable ultimo_error        : integer := 0;
    begin
        if (reloj'event and reloj='1') then
            contador := contador + 1;
            if (contador = 1000000) then -- Cada 10 ms => dt := 10/1000
                contador := 0;
                
                x_gyro_integer  := to_integer(signed( x_gyro ));
                y_gyro_integer  := to_integer(signed( y_gyro )) * 4;
                y_accel_integer := to_integer(signed( y_accel ));
                z_accel_integer := to_integer(signed( z_accel ));

                -- ``````````````````
                -- Filtrado
                angulo_crudo    := calc_angulo_crudo(y_accel_integer, z_accel_integer); -- atan ya está x1000;
                omega_dt        := (x_gyro_integer * decimales * dt / decimales) / gyro_gain; -- x_gyro / gyro_gain * dt
                angulo_filtrado := (A * (angulo_filtrado + omega_dt) + (decimales - A) * angulo_crudo) / decimales;

                -- ``````````````````
                -- PID
                error           := angulo_filtrado;                            -- Proporción
                sum_error       := sum_error + error * (dt / decimales);       -- Integración
                dErr            := (error - ultimo_error) / (dt / decimales);  -- Derivación
                velocidad       := (Kp * error + Ki * sum_error + Kd * dErr) / 100;
                ultimo_error    := error;
                
                velocidad_fin := velocidad / decimales;
                
                velocidad_a_temp := velocidad_fin - y_gyro_integer;
                velocidad_b_temp := velocidad_fin + y_gyro_integer;
                
                -- Evitar que la velocidad sobrepase el límite para PWM [0 - 255] con signo;
                if velocidad_a_temp > 255 then
                    velocidad_a_temp := 255;
                elsif velocidad_a_temp < -255 then
                    velocidad_a_temp := -255;
                end if;
                if velocidad_b_temp > 255 then
                    velocidad_b_temp := 255;
                elsif velocidad_b_temp < -255 then
                    velocidad_b_temp := -255;
                end if;
                
                velocidad_a_integer <= velocidad_a_temp;
                velocidad_b_integer <= velocidad_b_temp;

            end if;
        end if;
    end process;
    
    ajustar_Ks: process(reloj)
        variable Kp_ultimo_estado : std_logic := '0';
        variable Kd_ultimo_estado : std_logic := '0';
        variable Ki_ultimo_estado : std_logic := '0';
    begin
        if (reloj'event and reloj='1') then
            if(kpUp = '1' and Kp_ultimo_estado = '0') then
                KP <= KP + 10;
            end if;
            Kp_ultimo_estado := kpUp;
            if(kdUp = '1' and Kd_ultimo_estado = '0') then
                Kd <= Kd + 10;
            end if;
            Kd_ultimo_estado := kdUp;
            if(kiUp = '1' and Ki_ultimo_estado = '0') then
                Ki <= Ki + 1;
            end if;
            Ki_ultimo_estado := kiUp;
        end if;
    end process ajustar_Ks;

    -- Transformar velocidad de motores a PWM [0 - 255]
    velocidad_a <= std_logic_vector(to_unsigned(abs( velocidad_a_integer ), velocidad_a'length));
    velocidad_b <= std_logic_vector(to_unsigned(abs( velocidad_b_integer ), velocidad_b'length));
    
    -- Asignar el sentido de los motores para el puente H
    l298n_in1 <= '0' when velocidad_a_integer > 0 else '1';
    l298n_in2 <= '1' when velocidad_a_integer > 0 else '0';
    l298n_in3 <= '0' when velocidad_b_integer > 0 else '1';
    l298n_in4 <= '1' when velocidad_b_integer > 0 else '0';

end comportamiento;