

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity control_motores is
    Port ();

end control_motores;

architecture Comportamiento of decodificador_mpu6050 is

    
begin
    process(reloj)
    begin
        if (reloj'event and reloj='1') then

        end if;
    end process;
end Comportamiento;